
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h5b4f5272;
    ram_cell[       1] = 32'h0;  // 32'h31e36771;
    ram_cell[       2] = 32'h0;  // 32'h0630ac71;
    ram_cell[       3] = 32'h0;  // 32'h1253f8e2;
    ram_cell[       4] = 32'h0;  // 32'hb5763d64;
    ram_cell[       5] = 32'h0;  // 32'h7c582089;
    ram_cell[       6] = 32'h0;  // 32'hf3fac14e;
    ram_cell[       7] = 32'h0;  // 32'ha4aed99a;
    ram_cell[       8] = 32'h0;  // 32'h438d834e;
    ram_cell[       9] = 32'h0;  // 32'hf4584225;
    ram_cell[      10] = 32'h0;  // 32'hd883c1e6;
    ram_cell[      11] = 32'h0;  // 32'h04cefdd6;
    ram_cell[      12] = 32'h0;  // 32'hde41f82d;
    ram_cell[      13] = 32'h0;  // 32'h6057512b;
    ram_cell[      14] = 32'h0;  // 32'hf0d513c0;
    ram_cell[      15] = 32'h0;  // 32'h3282e7cf;
    ram_cell[      16] = 32'h0;  // 32'h51e716de;
    ram_cell[      17] = 32'h0;  // 32'h697d0ce8;
    ram_cell[      18] = 32'h0;  // 32'hfe90f66e;
    ram_cell[      19] = 32'h0;  // 32'h9d5bf4b7;
    ram_cell[      20] = 32'h0;  // 32'hdeec06fe;
    ram_cell[      21] = 32'h0;  // 32'h71c05274;
    ram_cell[      22] = 32'h0;  // 32'hf857745d;
    ram_cell[      23] = 32'h0;  // 32'hc90ba80f;
    ram_cell[      24] = 32'h0;  // 32'he74c52e0;
    ram_cell[      25] = 32'h0;  // 32'h59c04509;
    ram_cell[      26] = 32'h0;  // 32'he1814b45;
    ram_cell[      27] = 32'h0;  // 32'h336e30c8;
    ram_cell[      28] = 32'h0;  // 32'h615a10eb;
    ram_cell[      29] = 32'h0;  // 32'hea4119d8;
    ram_cell[      30] = 32'h0;  // 32'h8323691b;
    ram_cell[      31] = 32'h0;  // 32'h3eb60b2c;
    ram_cell[      32] = 32'h0;  // 32'h08b0b5b2;
    ram_cell[      33] = 32'h0;  // 32'h33f5cb69;
    ram_cell[      34] = 32'h0;  // 32'h37da30bc;
    ram_cell[      35] = 32'h0;  // 32'h4c28ec22;
    ram_cell[      36] = 32'h0;  // 32'hb6ba0ce0;
    ram_cell[      37] = 32'h0;  // 32'h38f53b88;
    ram_cell[      38] = 32'h0;  // 32'h4af82d15;
    ram_cell[      39] = 32'h0;  // 32'hd0622d41;
    ram_cell[      40] = 32'h0;  // 32'hf1a952a6;
    ram_cell[      41] = 32'h0;  // 32'hccac2be6;
    ram_cell[      42] = 32'h0;  // 32'h443aac0f;
    ram_cell[      43] = 32'h0;  // 32'h0a2e506a;
    ram_cell[      44] = 32'h0;  // 32'h9d18c129;
    ram_cell[      45] = 32'h0;  // 32'h7c533135;
    ram_cell[      46] = 32'h0;  // 32'h27f535d3;
    ram_cell[      47] = 32'h0;  // 32'h80b7eab3;
    ram_cell[      48] = 32'h0;  // 32'hdc353acb;
    ram_cell[      49] = 32'h0;  // 32'heb4f64cc;
    ram_cell[      50] = 32'h0;  // 32'h37df8bbc;
    ram_cell[      51] = 32'h0;  // 32'hd6eda759;
    ram_cell[      52] = 32'h0;  // 32'h009b3855;
    ram_cell[      53] = 32'h0;  // 32'h2b154c18;
    ram_cell[      54] = 32'h0;  // 32'h89c3cef5;
    ram_cell[      55] = 32'h0;  // 32'ha2c4559f;
    ram_cell[      56] = 32'h0;  // 32'h6e9a9ae5;
    ram_cell[      57] = 32'h0;  // 32'ha9541ad6;
    ram_cell[      58] = 32'h0;  // 32'h613a713e;
    ram_cell[      59] = 32'h0;  // 32'h99a3fc8b;
    ram_cell[      60] = 32'h0;  // 32'he7ed8938;
    ram_cell[      61] = 32'h0;  // 32'h5aedff61;
    ram_cell[      62] = 32'h0;  // 32'h97dc79d1;
    ram_cell[      63] = 32'h0;  // 32'he796eeb5;
    ram_cell[      64] = 32'h0;  // 32'h7e8f8e24;
    ram_cell[      65] = 32'h0;  // 32'ha3694631;
    ram_cell[      66] = 32'h0;  // 32'h3dc2f90b;
    ram_cell[      67] = 32'h0;  // 32'hc2274d8b;
    ram_cell[      68] = 32'h0;  // 32'ha599706a;
    ram_cell[      69] = 32'h0;  // 32'h2e777ef3;
    ram_cell[      70] = 32'h0;  // 32'hc991c22c;
    ram_cell[      71] = 32'h0;  // 32'h12c19303;
    ram_cell[      72] = 32'h0;  // 32'h5f5dec08;
    ram_cell[      73] = 32'h0;  // 32'he1bf5d38;
    ram_cell[      74] = 32'h0;  // 32'ha396b916;
    ram_cell[      75] = 32'h0;  // 32'hdd1257b3;
    ram_cell[      76] = 32'h0;  // 32'hd18a1913;
    ram_cell[      77] = 32'h0;  // 32'hb8858060;
    ram_cell[      78] = 32'h0;  // 32'h94fce898;
    ram_cell[      79] = 32'h0;  // 32'h18f6f6c7;
    ram_cell[      80] = 32'h0;  // 32'hf6d69347;
    ram_cell[      81] = 32'h0;  // 32'h001c4ca6;
    ram_cell[      82] = 32'h0;  // 32'h50e0a680;
    ram_cell[      83] = 32'h0;  // 32'h933addf5;
    ram_cell[      84] = 32'h0;  // 32'hc1b17fd1;
    ram_cell[      85] = 32'h0;  // 32'h6d8a0b9e;
    ram_cell[      86] = 32'h0;  // 32'hc47a0fe0;
    ram_cell[      87] = 32'h0;  // 32'h574a44b3;
    ram_cell[      88] = 32'h0;  // 32'h43b0f371;
    ram_cell[      89] = 32'h0;  // 32'hd2703668;
    ram_cell[      90] = 32'h0;  // 32'hf53105a0;
    ram_cell[      91] = 32'h0;  // 32'hc3f9fe00;
    ram_cell[      92] = 32'h0;  // 32'h91bcd20e;
    ram_cell[      93] = 32'h0;  // 32'ha2c1af13;
    ram_cell[      94] = 32'h0;  // 32'h40e6cf53;
    ram_cell[      95] = 32'h0;  // 32'hcc33485f;
    ram_cell[      96] = 32'h0;  // 32'hfff20c8e;
    ram_cell[      97] = 32'h0;  // 32'h19c4cd11;
    ram_cell[      98] = 32'h0;  // 32'h22ca98f5;
    ram_cell[      99] = 32'h0;  // 32'hd38e3e6d;
    ram_cell[     100] = 32'h0;  // 32'hf2aa8672;
    ram_cell[     101] = 32'h0;  // 32'h988f26f6;
    ram_cell[     102] = 32'h0;  // 32'h54c64f6a;
    ram_cell[     103] = 32'h0;  // 32'hd75741cb;
    ram_cell[     104] = 32'h0;  // 32'h14c8e87d;
    ram_cell[     105] = 32'h0;  // 32'h5e909e96;
    ram_cell[     106] = 32'h0;  // 32'h652640c5;
    ram_cell[     107] = 32'h0;  // 32'h29c9ef25;
    ram_cell[     108] = 32'h0;  // 32'hfc1470db;
    ram_cell[     109] = 32'h0;  // 32'h557f0b40;
    ram_cell[     110] = 32'h0;  // 32'he0412ed1;
    ram_cell[     111] = 32'h0;  // 32'h075b2178;
    ram_cell[     112] = 32'h0;  // 32'hbcc1f84b;
    ram_cell[     113] = 32'h0;  // 32'hf896a64f;
    ram_cell[     114] = 32'h0;  // 32'he4422eae;
    ram_cell[     115] = 32'h0;  // 32'he95b1d5d;
    ram_cell[     116] = 32'h0;  // 32'he524f48b;
    ram_cell[     117] = 32'h0;  // 32'h9313f39e;
    ram_cell[     118] = 32'h0;  // 32'h248170b1;
    ram_cell[     119] = 32'h0;  // 32'hc5cb20b5;
    ram_cell[     120] = 32'h0;  // 32'h408ea02b;
    ram_cell[     121] = 32'h0;  // 32'h5ac777d0;
    ram_cell[     122] = 32'h0;  // 32'ha064234e;
    ram_cell[     123] = 32'h0;  // 32'hcf6628b0;
    ram_cell[     124] = 32'h0;  // 32'h6f25919c;
    ram_cell[     125] = 32'h0;  // 32'h79820324;
    ram_cell[     126] = 32'h0;  // 32'h02b7132e;
    ram_cell[     127] = 32'h0;  // 32'h3bac1463;
    ram_cell[     128] = 32'h0;  // 32'ha8fc8608;
    ram_cell[     129] = 32'h0;  // 32'he0febae5;
    ram_cell[     130] = 32'h0;  // 32'h99074dbb;
    ram_cell[     131] = 32'h0;  // 32'ha0994b80;
    ram_cell[     132] = 32'h0;  // 32'heed06515;
    ram_cell[     133] = 32'h0;  // 32'h2fbe1180;
    ram_cell[     134] = 32'h0;  // 32'hfe685ced;
    ram_cell[     135] = 32'h0;  // 32'h2d1f060f;
    ram_cell[     136] = 32'h0;  // 32'hcc225275;
    ram_cell[     137] = 32'h0;  // 32'h87fce5bb;
    ram_cell[     138] = 32'h0;  // 32'h27d93327;
    ram_cell[     139] = 32'h0;  // 32'h1a37ba19;
    ram_cell[     140] = 32'h0;  // 32'hcb64a578;
    ram_cell[     141] = 32'h0;  // 32'h667db85a;
    ram_cell[     142] = 32'h0;  // 32'h4478afff;
    ram_cell[     143] = 32'h0;  // 32'h6b348382;
    ram_cell[     144] = 32'h0;  // 32'h4a391505;
    ram_cell[     145] = 32'h0;  // 32'habf77938;
    ram_cell[     146] = 32'h0;  // 32'h6231786d;
    ram_cell[     147] = 32'h0;  // 32'ha2a43905;
    ram_cell[     148] = 32'h0;  // 32'h10d7c55c;
    ram_cell[     149] = 32'h0;  // 32'h06a2f29a;
    ram_cell[     150] = 32'h0;  // 32'hc1169903;
    ram_cell[     151] = 32'h0;  // 32'h39ac9f67;
    ram_cell[     152] = 32'h0;  // 32'h24a056ad;
    ram_cell[     153] = 32'h0;  // 32'hbec18809;
    ram_cell[     154] = 32'h0;  // 32'hdbcd330c;
    ram_cell[     155] = 32'h0;  // 32'h2cd3807d;
    ram_cell[     156] = 32'h0;  // 32'h43966f4f;
    ram_cell[     157] = 32'h0;  // 32'hd3e16645;
    ram_cell[     158] = 32'h0;  // 32'he2a55eb6;
    ram_cell[     159] = 32'h0;  // 32'h30cd6515;
    ram_cell[     160] = 32'h0;  // 32'h8b3000f9;
    ram_cell[     161] = 32'h0;  // 32'h5048a8b4;
    ram_cell[     162] = 32'h0;  // 32'hfb007b41;
    ram_cell[     163] = 32'h0;  // 32'he0a51ce6;
    ram_cell[     164] = 32'h0;  // 32'h531feeea;
    ram_cell[     165] = 32'h0;  // 32'hd9432b9d;
    ram_cell[     166] = 32'h0;  // 32'h01901247;
    ram_cell[     167] = 32'h0;  // 32'hb97b65e9;
    ram_cell[     168] = 32'h0;  // 32'hcd0047db;
    ram_cell[     169] = 32'h0;  // 32'h86dc02b4;
    ram_cell[     170] = 32'h0;  // 32'h38333f4b;
    ram_cell[     171] = 32'h0;  // 32'hb1b29dc4;
    ram_cell[     172] = 32'h0;  // 32'hc0fffdce;
    ram_cell[     173] = 32'h0;  // 32'he1dac616;
    ram_cell[     174] = 32'h0;  // 32'h746da07e;
    ram_cell[     175] = 32'h0;  // 32'h11e3a981;
    ram_cell[     176] = 32'h0;  // 32'h2651a5f0;
    ram_cell[     177] = 32'h0;  // 32'h0582ffde;
    ram_cell[     178] = 32'h0;  // 32'h00acb7f0;
    ram_cell[     179] = 32'h0;  // 32'hf3ae5c15;
    ram_cell[     180] = 32'h0;  // 32'h05db1b1c;
    ram_cell[     181] = 32'h0;  // 32'h136e6dfd;
    ram_cell[     182] = 32'h0;  // 32'he1728505;
    ram_cell[     183] = 32'h0;  // 32'h4d42c89d;
    ram_cell[     184] = 32'h0;  // 32'ha1b814fe;
    ram_cell[     185] = 32'h0;  // 32'hb72d6870;
    ram_cell[     186] = 32'h0;  // 32'hf62ecabe;
    ram_cell[     187] = 32'h0;  // 32'hb481e39c;
    ram_cell[     188] = 32'h0;  // 32'hd2d0f70c;
    ram_cell[     189] = 32'h0;  // 32'hf55eaa8f;
    ram_cell[     190] = 32'h0;  // 32'h2cdac20c;
    ram_cell[     191] = 32'h0;  // 32'h927a7e62;
    ram_cell[     192] = 32'h0;  // 32'h35e14e27;
    ram_cell[     193] = 32'h0;  // 32'h4e1cbd22;
    ram_cell[     194] = 32'h0;  // 32'h77e87143;
    ram_cell[     195] = 32'h0;  // 32'h2b823444;
    ram_cell[     196] = 32'h0;  // 32'h3bd4dbeb;
    ram_cell[     197] = 32'h0;  // 32'hae27b6fc;
    ram_cell[     198] = 32'h0;  // 32'h3e06fb56;
    ram_cell[     199] = 32'h0;  // 32'h80b73f99;
    ram_cell[     200] = 32'h0;  // 32'h863acb6b;
    ram_cell[     201] = 32'h0;  // 32'he9c1926a;
    ram_cell[     202] = 32'h0;  // 32'h928fca80;
    ram_cell[     203] = 32'h0;  // 32'h84167d40;
    ram_cell[     204] = 32'h0;  // 32'h4810313c;
    ram_cell[     205] = 32'h0;  // 32'h1a078945;
    ram_cell[     206] = 32'h0;  // 32'h5624da5d;
    ram_cell[     207] = 32'h0;  // 32'hd9cfd208;
    ram_cell[     208] = 32'h0;  // 32'hffc6601f;
    ram_cell[     209] = 32'h0;  // 32'h701d7b2d;
    ram_cell[     210] = 32'h0;  // 32'ha5aec90d;
    ram_cell[     211] = 32'h0;  // 32'h517b6459;
    ram_cell[     212] = 32'h0;  // 32'h2b546413;
    ram_cell[     213] = 32'h0;  // 32'h1f4adfbd;
    ram_cell[     214] = 32'h0;  // 32'h5cf7cd7d;
    ram_cell[     215] = 32'h0;  // 32'ha46b0579;
    ram_cell[     216] = 32'h0;  // 32'h77957992;
    ram_cell[     217] = 32'h0;  // 32'h4eef7998;
    ram_cell[     218] = 32'h0;  // 32'hfd63c2d8;
    ram_cell[     219] = 32'h0;  // 32'h555f0328;
    ram_cell[     220] = 32'h0;  // 32'h2dc9fc29;
    ram_cell[     221] = 32'h0;  // 32'hae489606;
    ram_cell[     222] = 32'h0;  // 32'ha5613660;
    ram_cell[     223] = 32'h0;  // 32'h9194ab53;
    ram_cell[     224] = 32'h0;  // 32'h735bb971;
    ram_cell[     225] = 32'h0;  // 32'hdbe5fdfd;
    ram_cell[     226] = 32'h0;  // 32'he9a7b4bb;
    ram_cell[     227] = 32'h0;  // 32'h65ea1b75;
    ram_cell[     228] = 32'h0;  // 32'ha25671fd;
    ram_cell[     229] = 32'h0;  // 32'hebc0c460;
    ram_cell[     230] = 32'h0;  // 32'he7b23b20;
    ram_cell[     231] = 32'h0;  // 32'h56762b46;
    ram_cell[     232] = 32'h0;  // 32'hc985d7be;
    ram_cell[     233] = 32'h0;  // 32'hf5172315;
    ram_cell[     234] = 32'h0;  // 32'ha97b095e;
    ram_cell[     235] = 32'h0;  // 32'h284568a7;
    ram_cell[     236] = 32'h0;  // 32'h1b95160f;
    ram_cell[     237] = 32'h0;  // 32'h0b4f7bd4;
    ram_cell[     238] = 32'h0;  // 32'hec89c1d9;
    ram_cell[     239] = 32'h0;  // 32'he50652d1;
    ram_cell[     240] = 32'h0;  // 32'he0e28ba5;
    ram_cell[     241] = 32'h0;  // 32'hc3dc9a45;
    ram_cell[     242] = 32'h0;  // 32'he87031c7;
    ram_cell[     243] = 32'h0;  // 32'h668b0bb9;
    ram_cell[     244] = 32'h0;  // 32'h79d8cfd3;
    ram_cell[     245] = 32'h0;  // 32'hb038a5c7;
    ram_cell[     246] = 32'h0;  // 32'h471a7b76;
    ram_cell[     247] = 32'h0;  // 32'he4b5c4e4;
    ram_cell[     248] = 32'h0;  // 32'h2b7cbd3b;
    ram_cell[     249] = 32'h0;  // 32'h6e7bd705;
    ram_cell[     250] = 32'h0;  // 32'h6e72e622;
    ram_cell[     251] = 32'h0;  // 32'h3381ed93;
    ram_cell[     252] = 32'h0;  // 32'h750de595;
    ram_cell[     253] = 32'h0;  // 32'h79ae2214;
    ram_cell[     254] = 32'h0;  // 32'h85cf7e49;
    ram_cell[     255] = 32'h0;  // 32'h5952717b;
    // src matrix A
    ram_cell[     256] = 32'hf3f08ab9;
    ram_cell[     257] = 32'h069ac97a;
    ram_cell[     258] = 32'h3b5dd9bc;
    ram_cell[     259] = 32'h43e0836f;
    ram_cell[     260] = 32'h3b971806;
    ram_cell[     261] = 32'ha3895853;
    ram_cell[     262] = 32'hc053509e;
    ram_cell[     263] = 32'h3a865575;
    ram_cell[     264] = 32'h5e10f84e;
    ram_cell[     265] = 32'h0f486db3;
    ram_cell[     266] = 32'h2b492017;
    ram_cell[     267] = 32'hdef437ad;
    ram_cell[     268] = 32'h3c6b89c8;
    ram_cell[     269] = 32'hcdea939e;
    ram_cell[     270] = 32'hcd5bef97;
    ram_cell[     271] = 32'hf55a2a25;
    ram_cell[     272] = 32'h667bff57;
    ram_cell[     273] = 32'h8de9d679;
    ram_cell[     274] = 32'h78218fd5;
    ram_cell[     275] = 32'h08df8fa2;
    ram_cell[     276] = 32'h6be41ef2;
    ram_cell[     277] = 32'h37252116;
    ram_cell[     278] = 32'h8bea8ad1;
    ram_cell[     279] = 32'he35d4a4a;
    ram_cell[     280] = 32'hf4262ad8;
    ram_cell[     281] = 32'h65a04117;
    ram_cell[     282] = 32'h6a56d3f0;
    ram_cell[     283] = 32'hfe310e24;
    ram_cell[     284] = 32'hfcdd65d6;
    ram_cell[     285] = 32'h0108b563;
    ram_cell[     286] = 32'hbdaa7f66;
    ram_cell[     287] = 32'h8ef16159;
    ram_cell[     288] = 32'hce424acf;
    ram_cell[     289] = 32'h13373979;
    ram_cell[     290] = 32'h6c2f9c55;
    ram_cell[     291] = 32'h1d8e6828;
    ram_cell[     292] = 32'ha2106fe9;
    ram_cell[     293] = 32'h6736e50d;
    ram_cell[     294] = 32'hb546953e;
    ram_cell[     295] = 32'hccd3acdf;
    ram_cell[     296] = 32'hcb2ee877;
    ram_cell[     297] = 32'hf0139b34;
    ram_cell[     298] = 32'h7c48e3b0;
    ram_cell[     299] = 32'haf5be650;
    ram_cell[     300] = 32'h5452d04a;
    ram_cell[     301] = 32'h5f374e7c;
    ram_cell[     302] = 32'h64a3815b;
    ram_cell[     303] = 32'hfe2c5bb5;
    ram_cell[     304] = 32'h411fadee;
    ram_cell[     305] = 32'h49b296d7;
    ram_cell[     306] = 32'hb7ac32ca;
    ram_cell[     307] = 32'h626a37b2;
    ram_cell[     308] = 32'h982fc174;
    ram_cell[     309] = 32'h545f7863;
    ram_cell[     310] = 32'h3bb5d248;
    ram_cell[     311] = 32'h87b200b3;
    ram_cell[     312] = 32'hacf8b065;
    ram_cell[     313] = 32'h0ec95bdb;
    ram_cell[     314] = 32'h20bbafb8;
    ram_cell[     315] = 32'hc1f7abe0;
    ram_cell[     316] = 32'h1a104702;
    ram_cell[     317] = 32'h32937c8b;
    ram_cell[     318] = 32'h2b7e9dce;
    ram_cell[     319] = 32'h2455afa1;
    ram_cell[     320] = 32'hd99eafef;
    ram_cell[     321] = 32'hfd5e2fab;
    ram_cell[     322] = 32'hffe106bb;
    ram_cell[     323] = 32'h7c9e9a6d;
    ram_cell[     324] = 32'h159f4e12;
    ram_cell[     325] = 32'h9cecb46d;
    ram_cell[     326] = 32'h4154642d;
    ram_cell[     327] = 32'hc29b7806;
    ram_cell[     328] = 32'h95628aaa;
    ram_cell[     329] = 32'h75e2b461;
    ram_cell[     330] = 32'h8e27ca8d;
    ram_cell[     331] = 32'h7c885e58;
    ram_cell[     332] = 32'hf285bbb5;
    ram_cell[     333] = 32'hee882e78;
    ram_cell[     334] = 32'h13355f33;
    ram_cell[     335] = 32'h8d0fbcf2;
    ram_cell[     336] = 32'he8965d03;
    ram_cell[     337] = 32'h7c6c5ab3;
    ram_cell[     338] = 32'h4180a1ee;
    ram_cell[     339] = 32'hf5d7d2ba;
    ram_cell[     340] = 32'hf8a8d6e0;
    ram_cell[     341] = 32'h21045bc7;
    ram_cell[     342] = 32'h86319953;
    ram_cell[     343] = 32'ha4ea8bdf;
    ram_cell[     344] = 32'h43002135;
    ram_cell[     345] = 32'h11d50e54;
    ram_cell[     346] = 32'h3e41bfe4;
    ram_cell[     347] = 32'h605c17ca;
    ram_cell[     348] = 32'hce0e746e;
    ram_cell[     349] = 32'hb9865d9b;
    ram_cell[     350] = 32'h72c7e1cc;
    ram_cell[     351] = 32'hb945cbc2;
    ram_cell[     352] = 32'haa5a0705;
    ram_cell[     353] = 32'h72706a78;
    ram_cell[     354] = 32'he7c0638c;
    ram_cell[     355] = 32'h1db924b6;
    ram_cell[     356] = 32'h44e6b175;
    ram_cell[     357] = 32'hdc1afb3a;
    ram_cell[     358] = 32'h63c82ada;
    ram_cell[     359] = 32'h96b120a6;
    ram_cell[     360] = 32'h4823ebf5;
    ram_cell[     361] = 32'h03216cef;
    ram_cell[     362] = 32'h8e213a3a;
    ram_cell[     363] = 32'h64ade210;
    ram_cell[     364] = 32'h140e7250;
    ram_cell[     365] = 32'h09443224;
    ram_cell[     366] = 32'hc62f11d4;
    ram_cell[     367] = 32'h2fe7ab9a;
    ram_cell[     368] = 32'he9bef4d2;
    ram_cell[     369] = 32'h9200cb24;
    ram_cell[     370] = 32'h38438ebd;
    ram_cell[     371] = 32'h8c3af9f1;
    ram_cell[     372] = 32'hbdf4372d;
    ram_cell[     373] = 32'hf3f6d336;
    ram_cell[     374] = 32'h3349b858;
    ram_cell[     375] = 32'h4bf584a2;
    ram_cell[     376] = 32'h526365af;
    ram_cell[     377] = 32'h99215da4;
    ram_cell[     378] = 32'h893e0ac1;
    ram_cell[     379] = 32'h93d82780;
    ram_cell[     380] = 32'h0876b404;
    ram_cell[     381] = 32'h0c54ecf4;
    ram_cell[     382] = 32'ha6a1ac68;
    ram_cell[     383] = 32'hacd26017;
    ram_cell[     384] = 32'h3817c0b4;
    ram_cell[     385] = 32'h66bf0b00;
    ram_cell[     386] = 32'hb7e3ed40;
    ram_cell[     387] = 32'h18932f63;
    ram_cell[     388] = 32'h361da84a;
    ram_cell[     389] = 32'hccff9bdf;
    ram_cell[     390] = 32'h94646bc6;
    ram_cell[     391] = 32'hbd3aa227;
    ram_cell[     392] = 32'hc575adbd;
    ram_cell[     393] = 32'h67fb726b;
    ram_cell[     394] = 32'h8d05639f;
    ram_cell[     395] = 32'h388b47de;
    ram_cell[     396] = 32'h9ee675cf;
    ram_cell[     397] = 32'h2026ab88;
    ram_cell[     398] = 32'hd0ac07b3;
    ram_cell[     399] = 32'h78bd26d2;
    ram_cell[     400] = 32'h8cfabb45;
    ram_cell[     401] = 32'h73678bac;
    ram_cell[     402] = 32'h90da5245;
    ram_cell[     403] = 32'hc88783a0;
    ram_cell[     404] = 32'h20f0e48e;
    ram_cell[     405] = 32'ha1aa2d78;
    ram_cell[     406] = 32'h8d85a422;
    ram_cell[     407] = 32'h69bfb502;
    ram_cell[     408] = 32'h2290e9fd;
    ram_cell[     409] = 32'hb381f53e;
    ram_cell[     410] = 32'h7039e51f;
    ram_cell[     411] = 32'ha6519851;
    ram_cell[     412] = 32'hb2c455b0;
    ram_cell[     413] = 32'hc062e72d;
    ram_cell[     414] = 32'h95814ee2;
    ram_cell[     415] = 32'hc90c9ef5;
    ram_cell[     416] = 32'h1c11156d;
    ram_cell[     417] = 32'hc1ba86d0;
    ram_cell[     418] = 32'h406b0337;
    ram_cell[     419] = 32'h165a0e51;
    ram_cell[     420] = 32'h94d01baa;
    ram_cell[     421] = 32'h259378e0;
    ram_cell[     422] = 32'hdd98d8f5;
    ram_cell[     423] = 32'h0268cec4;
    ram_cell[     424] = 32'h7cf2b8ab;
    ram_cell[     425] = 32'h6759da63;
    ram_cell[     426] = 32'hb6a96050;
    ram_cell[     427] = 32'h636a73f8;
    ram_cell[     428] = 32'h1e3f3175;
    ram_cell[     429] = 32'h891ba716;
    ram_cell[     430] = 32'h4c5358f3;
    ram_cell[     431] = 32'h7ad1a9ae;
    ram_cell[     432] = 32'hc526f4b6;
    ram_cell[     433] = 32'h7d6ae84e;
    ram_cell[     434] = 32'hf2f2769e;
    ram_cell[     435] = 32'hf5c68534;
    ram_cell[     436] = 32'h9d0fbc09;
    ram_cell[     437] = 32'hbb4d338b;
    ram_cell[     438] = 32'haedfb076;
    ram_cell[     439] = 32'h31cf35f0;
    ram_cell[     440] = 32'h711e0fc2;
    ram_cell[     441] = 32'h8dbffe56;
    ram_cell[     442] = 32'h16bf05b1;
    ram_cell[     443] = 32'hcb0ddb37;
    ram_cell[     444] = 32'h6b26a907;
    ram_cell[     445] = 32'hf44a6f15;
    ram_cell[     446] = 32'h7ff7ef8d;
    ram_cell[     447] = 32'hc3057ae7;
    ram_cell[     448] = 32'h4d52cd67;
    ram_cell[     449] = 32'hf027a76d;
    ram_cell[     450] = 32'h9c217537;
    ram_cell[     451] = 32'h6b458bb9;
    ram_cell[     452] = 32'h5cd67eae;
    ram_cell[     453] = 32'h2e6cfb48;
    ram_cell[     454] = 32'h212a36f1;
    ram_cell[     455] = 32'h5a9439aa;
    ram_cell[     456] = 32'h2cb41ac9;
    ram_cell[     457] = 32'hef88e071;
    ram_cell[     458] = 32'ha18e103a;
    ram_cell[     459] = 32'hb6ea030d;
    ram_cell[     460] = 32'h72419378;
    ram_cell[     461] = 32'h53f815ca;
    ram_cell[     462] = 32'h4cc8650d;
    ram_cell[     463] = 32'h58972435;
    ram_cell[     464] = 32'hc9ca3a88;
    ram_cell[     465] = 32'h2289c333;
    ram_cell[     466] = 32'h4ceac55d;
    ram_cell[     467] = 32'h8a27c758;
    ram_cell[     468] = 32'h818a564c;
    ram_cell[     469] = 32'h018e9399;
    ram_cell[     470] = 32'ha6649910;
    ram_cell[     471] = 32'h8fd7fe12;
    ram_cell[     472] = 32'h5dfd1aae;
    ram_cell[     473] = 32'h4248b9de;
    ram_cell[     474] = 32'h3b450c43;
    ram_cell[     475] = 32'hb37f0d75;
    ram_cell[     476] = 32'h28e818ca;
    ram_cell[     477] = 32'h59379f67;
    ram_cell[     478] = 32'h78a5b6dc;
    ram_cell[     479] = 32'hf274fd39;
    ram_cell[     480] = 32'hf0d397d2;
    ram_cell[     481] = 32'h7f9a6cac;
    ram_cell[     482] = 32'h00e5444b;
    ram_cell[     483] = 32'h75c7df51;
    ram_cell[     484] = 32'h09f1e54b;
    ram_cell[     485] = 32'hd5e696c1;
    ram_cell[     486] = 32'h4838f1ba;
    ram_cell[     487] = 32'h41685ce9;
    ram_cell[     488] = 32'hffab8d45;
    ram_cell[     489] = 32'h81b7c1c4;
    ram_cell[     490] = 32'hb9d7334e;
    ram_cell[     491] = 32'h12be4ed9;
    ram_cell[     492] = 32'hcfaad3ac;
    ram_cell[     493] = 32'hedae7847;
    ram_cell[     494] = 32'h5927789c;
    ram_cell[     495] = 32'hb0b969e3;
    ram_cell[     496] = 32'hfaebc5d1;
    ram_cell[     497] = 32'hbab1a876;
    ram_cell[     498] = 32'h539159ff;
    ram_cell[     499] = 32'h7f011eda;
    ram_cell[     500] = 32'haa95c86d;
    ram_cell[     501] = 32'h28f47b4e;
    ram_cell[     502] = 32'h90adf519;
    ram_cell[     503] = 32'hf7debc0b;
    ram_cell[     504] = 32'h3a260bcc;
    ram_cell[     505] = 32'h951bdd44;
    ram_cell[     506] = 32'ha078a4ad;
    ram_cell[     507] = 32'h28239f35;
    ram_cell[     508] = 32'hdf619ebd;
    ram_cell[     509] = 32'h62fd718f;
    ram_cell[     510] = 32'h8636f878;
    ram_cell[     511] = 32'hb9dde5d9;
    // src matrix B
    ram_cell[     512] = 32'h8882d28f;
    ram_cell[     513] = 32'h46cf74a8;
    ram_cell[     514] = 32'ha601f279;
    ram_cell[     515] = 32'ha8ad5437;
    ram_cell[     516] = 32'h10526e61;
    ram_cell[     517] = 32'hd0ff495d;
    ram_cell[     518] = 32'h9014624e;
    ram_cell[     519] = 32'h71bc8c28;
    ram_cell[     520] = 32'h38b362ff;
    ram_cell[     521] = 32'h67e768d2;
    ram_cell[     522] = 32'h1c832152;
    ram_cell[     523] = 32'h8000d8f5;
    ram_cell[     524] = 32'h2da3848f;
    ram_cell[     525] = 32'h1abd55a3;
    ram_cell[     526] = 32'hedb57e2d;
    ram_cell[     527] = 32'h6106abf0;
    ram_cell[     528] = 32'hfb94855b;
    ram_cell[     529] = 32'h84475a01;
    ram_cell[     530] = 32'h6486ed3a;
    ram_cell[     531] = 32'h354db5df;
    ram_cell[     532] = 32'h39a590f1;
    ram_cell[     533] = 32'h01be32fe;
    ram_cell[     534] = 32'h70d7cd0f;
    ram_cell[     535] = 32'h7556074b;
    ram_cell[     536] = 32'h20bc1062;
    ram_cell[     537] = 32'h0ca1407d;
    ram_cell[     538] = 32'h407c9774;
    ram_cell[     539] = 32'h7ea918d7;
    ram_cell[     540] = 32'h7f62b105;
    ram_cell[     541] = 32'hcbe4213e;
    ram_cell[     542] = 32'h6e7696fd;
    ram_cell[     543] = 32'hbfe69e88;
    ram_cell[     544] = 32'hac5666fe;
    ram_cell[     545] = 32'h5d7658f7;
    ram_cell[     546] = 32'h4d6560d5;
    ram_cell[     547] = 32'heae86012;
    ram_cell[     548] = 32'h7de7377b;
    ram_cell[     549] = 32'h9d6d22bd;
    ram_cell[     550] = 32'h2d1ae58d;
    ram_cell[     551] = 32'h4fd632c9;
    ram_cell[     552] = 32'h9bf5d669;
    ram_cell[     553] = 32'h2243346c;
    ram_cell[     554] = 32'hb248cfda;
    ram_cell[     555] = 32'h99d6bb7f;
    ram_cell[     556] = 32'h0154a590;
    ram_cell[     557] = 32'h2a207635;
    ram_cell[     558] = 32'had95e9c6;
    ram_cell[     559] = 32'h53e10489;
    ram_cell[     560] = 32'hb80268d1;
    ram_cell[     561] = 32'head2f9a8;
    ram_cell[     562] = 32'hd0dccc49;
    ram_cell[     563] = 32'hd1fa07ee;
    ram_cell[     564] = 32'h97ca0eab;
    ram_cell[     565] = 32'hd19aaeda;
    ram_cell[     566] = 32'h350ad88d;
    ram_cell[     567] = 32'h38f70415;
    ram_cell[     568] = 32'h72723583;
    ram_cell[     569] = 32'he087f6b3;
    ram_cell[     570] = 32'hb620e135;
    ram_cell[     571] = 32'he9bf6fed;
    ram_cell[     572] = 32'h5f909182;
    ram_cell[     573] = 32'h2b2a12ad;
    ram_cell[     574] = 32'hc52c09bb;
    ram_cell[     575] = 32'h2f360bd0;
    ram_cell[     576] = 32'hb58f0362;
    ram_cell[     577] = 32'h2072a666;
    ram_cell[     578] = 32'h9a245c24;
    ram_cell[     579] = 32'hee69567e;
    ram_cell[     580] = 32'hc58b9807;
    ram_cell[     581] = 32'h2dc954a7;
    ram_cell[     582] = 32'h4b27be6a;
    ram_cell[     583] = 32'h00fee7d7;
    ram_cell[     584] = 32'hec2cce16;
    ram_cell[     585] = 32'he8dcd8e2;
    ram_cell[     586] = 32'hfcedfb74;
    ram_cell[     587] = 32'h0c5317bc;
    ram_cell[     588] = 32'h30d940c5;
    ram_cell[     589] = 32'h709fd433;
    ram_cell[     590] = 32'h7862a5da;
    ram_cell[     591] = 32'h071acad2;
    ram_cell[     592] = 32'ha191e892;
    ram_cell[     593] = 32'ha4e5c989;
    ram_cell[     594] = 32'h73438814;
    ram_cell[     595] = 32'hc2daf73e;
    ram_cell[     596] = 32'h66203f95;
    ram_cell[     597] = 32'h0ea8b787;
    ram_cell[     598] = 32'hd60a6296;
    ram_cell[     599] = 32'haa759ddf;
    ram_cell[     600] = 32'h26ee4a98;
    ram_cell[     601] = 32'h40d349cb;
    ram_cell[     602] = 32'h42f9a36c;
    ram_cell[     603] = 32'h0255d7a6;
    ram_cell[     604] = 32'ha71227cd;
    ram_cell[     605] = 32'h382398df;
    ram_cell[     606] = 32'h51636c0a;
    ram_cell[     607] = 32'h9d7362b6;
    ram_cell[     608] = 32'hdd89c69a;
    ram_cell[     609] = 32'h64d43585;
    ram_cell[     610] = 32'h5d0e24e0;
    ram_cell[     611] = 32'h9a5be40c;
    ram_cell[     612] = 32'hd74a8c01;
    ram_cell[     613] = 32'hac1cf059;
    ram_cell[     614] = 32'h155738d3;
    ram_cell[     615] = 32'h9898f7ae;
    ram_cell[     616] = 32'h75da6cfd;
    ram_cell[     617] = 32'h6a03a786;
    ram_cell[     618] = 32'h3f7280ab;
    ram_cell[     619] = 32'h693f7eff;
    ram_cell[     620] = 32'h1a353ec9;
    ram_cell[     621] = 32'h7bce50fc;
    ram_cell[     622] = 32'hc98ccb6f;
    ram_cell[     623] = 32'h3aca9d44;
    ram_cell[     624] = 32'hd69d116a;
    ram_cell[     625] = 32'he97d7e4e;
    ram_cell[     626] = 32'hbc52f0b5;
    ram_cell[     627] = 32'h5a554cff;
    ram_cell[     628] = 32'hbf476281;
    ram_cell[     629] = 32'h114b95c1;
    ram_cell[     630] = 32'h695553d5;
    ram_cell[     631] = 32'hb968de62;
    ram_cell[     632] = 32'he36f3b22;
    ram_cell[     633] = 32'h7ac59fad;
    ram_cell[     634] = 32'hf5582dd2;
    ram_cell[     635] = 32'h69e49191;
    ram_cell[     636] = 32'hd3e3fc9f;
    ram_cell[     637] = 32'h6af434cf;
    ram_cell[     638] = 32'hf135d240;
    ram_cell[     639] = 32'h718798ce;
    ram_cell[     640] = 32'h9a223860;
    ram_cell[     641] = 32'h1cf12fb5;
    ram_cell[     642] = 32'hf32920f3;
    ram_cell[     643] = 32'ha5ef3f62;
    ram_cell[     644] = 32'hca1eda9a;
    ram_cell[     645] = 32'h62863bbd;
    ram_cell[     646] = 32'h6d338f93;
    ram_cell[     647] = 32'h5b3e3272;
    ram_cell[     648] = 32'hd8f47a2e;
    ram_cell[     649] = 32'h98228bbf;
    ram_cell[     650] = 32'hfbc11788;
    ram_cell[     651] = 32'hd7f80b0f;
    ram_cell[     652] = 32'hd32941c1;
    ram_cell[     653] = 32'hc21fd16f;
    ram_cell[     654] = 32'hde33ce2c;
    ram_cell[     655] = 32'hed4b7168;
    ram_cell[     656] = 32'h3c0fdbe7;
    ram_cell[     657] = 32'ha3ba3b52;
    ram_cell[     658] = 32'h2d217f45;
    ram_cell[     659] = 32'h249acd30;
    ram_cell[     660] = 32'hf2ec6510;
    ram_cell[     661] = 32'h0ba3ea09;
    ram_cell[     662] = 32'h70adbeb9;
    ram_cell[     663] = 32'h96989dde;
    ram_cell[     664] = 32'hd05f1de4;
    ram_cell[     665] = 32'ha1748d43;
    ram_cell[     666] = 32'h2d25210d;
    ram_cell[     667] = 32'hf8050c97;
    ram_cell[     668] = 32'h6a1878d8;
    ram_cell[     669] = 32'ha6313b11;
    ram_cell[     670] = 32'h03ed827c;
    ram_cell[     671] = 32'h0cf0697c;
    ram_cell[     672] = 32'ha53eb0d0;
    ram_cell[     673] = 32'h7144527a;
    ram_cell[     674] = 32'h980fc18f;
    ram_cell[     675] = 32'hb5ee4782;
    ram_cell[     676] = 32'h6c2a3558;
    ram_cell[     677] = 32'hcc35d9ae;
    ram_cell[     678] = 32'h95ab3b67;
    ram_cell[     679] = 32'he6b82dd2;
    ram_cell[     680] = 32'h0e8aa2b7;
    ram_cell[     681] = 32'h51c650eb;
    ram_cell[     682] = 32'hc0957925;
    ram_cell[     683] = 32'h16bf6f15;
    ram_cell[     684] = 32'h2ad6437e;
    ram_cell[     685] = 32'hadc074cc;
    ram_cell[     686] = 32'hb05e4155;
    ram_cell[     687] = 32'h2aac5012;
    ram_cell[     688] = 32'hc0bea937;
    ram_cell[     689] = 32'h3509308f;
    ram_cell[     690] = 32'h42d090a2;
    ram_cell[     691] = 32'h0e20f6b5;
    ram_cell[     692] = 32'hbd7c0768;
    ram_cell[     693] = 32'hab64d69f;
    ram_cell[     694] = 32'h3193c45d;
    ram_cell[     695] = 32'h335e1fef;
    ram_cell[     696] = 32'h4f51fd9f;
    ram_cell[     697] = 32'h39d0bc68;
    ram_cell[     698] = 32'hcc0b69d6;
    ram_cell[     699] = 32'h63726498;
    ram_cell[     700] = 32'hca53a9b3;
    ram_cell[     701] = 32'h83636647;
    ram_cell[     702] = 32'h5e15b898;
    ram_cell[     703] = 32'hc7937319;
    ram_cell[     704] = 32'h5acfb050;
    ram_cell[     705] = 32'h92f54bef;
    ram_cell[     706] = 32'h9ca0c04c;
    ram_cell[     707] = 32'hb3497e29;
    ram_cell[     708] = 32'h076984d0;
    ram_cell[     709] = 32'h62506de5;
    ram_cell[     710] = 32'he9ca55f2;
    ram_cell[     711] = 32'hdb10d6b0;
    ram_cell[     712] = 32'h22cd4ae1;
    ram_cell[     713] = 32'h8c8cac38;
    ram_cell[     714] = 32'h1ee4ffff;
    ram_cell[     715] = 32'hb8c13109;
    ram_cell[     716] = 32'hdb004a9a;
    ram_cell[     717] = 32'h8dd33744;
    ram_cell[     718] = 32'h264a1312;
    ram_cell[     719] = 32'h70d12474;
    ram_cell[     720] = 32'h8cbec027;
    ram_cell[     721] = 32'h06e5ebc0;
    ram_cell[     722] = 32'hc75eaca1;
    ram_cell[     723] = 32'h1d8061aa;
    ram_cell[     724] = 32'h502200b2;
    ram_cell[     725] = 32'ha79ec8d9;
    ram_cell[     726] = 32'h91c3b880;
    ram_cell[     727] = 32'h9b858bbb;
    ram_cell[     728] = 32'h234048cb;
    ram_cell[     729] = 32'h9d501892;
    ram_cell[     730] = 32'he6a7fedf;
    ram_cell[     731] = 32'ha187eb7b;
    ram_cell[     732] = 32'heeffcf1c;
    ram_cell[     733] = 32'h3348068d;
    ram_cell[     734] = 32'had51026c;
    ram_cell[     735] = 32'hef719d91;
    ram_cell[     736] = 32'h1a69882e;
    ram_cell[     737] = 32'h3c608128;
    ram_cell[     738] = 32'ha1458e82;
    ram_cell[     739] = 32'h655c69fc;
    ram_cell[     740] = 32'h465a47b8;
    ram_cell[     741] = 32'h59dac69d;
    ram_cell[     742] = 32'h2ab57de8;
    ram_cell[     743] = 32'hc19b00c7;
    ram_cell[     744] = 32'h63b918fe;
    ram_cell[     745] = 32'hf6006d2f;
    ram_cell[     746] = 32'h16af46db;
    ram_cell[     747] = 32'hb0fd3715;
    ram_cell[     748] = 32'h95960f49;
    ram_cell[     749] = 32'h4cfe24a5;
    ram_cell[     750] = 32'h80c3da1d;
    ram_cell[     751] = 32'he9e4b0f0;
    ram_cell[     752] = 32'h55dc6928;
    ram_cell[     753] = 32'hf06a98ab;
    ram_cell[     754] = 32'h56bdc2e4;
    ram_cell[     755] = 32'h0890f1c9;
    ram_cell[     756] = 32'hb0bb563e;
    ram_cell[     757] = 32'hcffb5d91;
    ram_cell[     758] = 32'h748c376b;
    ram_cell[     759] = 32'hd3814da8;
    ram_cell[     760] = 32'hfefda04e;
    ram_cell[     761] = 32'hf705f39b;
    ram_cell[     762] = 32'h12b21750;
    ram_cell[     763] = 32'hdea1de90;
    ram_cell[     764] = 32'hd1113e16;
    ram_cell[     765] = 32'h17368980;
    ram_cell[     766] = 32'h6c7321a6;
    ram_cell[     767] = 32'hf089fb42;
end

endmodule

